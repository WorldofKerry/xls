module __adler32__add_two_f32(
  input wire clk,
  input wire [31:0] a,
  input wire [31:0] b,
  output wire [31:0] out
);
  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_a;
  reg [31:0] p0_b;
  always_ff @ (posedge clk) begin
    p0_a <= a;
    p0_b <= b;
  end

  // ===== Pipe stage 1:
  wire [7:0] p1_b_bexp__2_comb;
  wire [7:0] p1_a_bexp__2_comb;
  wire [8:0] p1_sum_comb;
  wire [22:0] p1_tuple_index_1463_comb;
  wire [22:0] p1_tuple_index_1464_comb;
  wire [7:0] p1_y_bexp_comb;
  wire [22:0] p1_y_fraction_comb;
  wire [7:0] p1_incremented_sum__1_comb;
  wire [27:0] p1_wide_y_comb;
  wire [7:0] p1_a_bexpbs_difference__1_comb;
  wire [7:0] p1_x_bexp_comb;
  wire [27:0] p1_wide_y__1_comb;
  wire [7:0] p1_sub_1482_comb;
  wire [22:0] p1_x_fraction_comb;
  wire [27:0] p1_dropped_comb;
  wire [27:0] p1_wide_x_comb;
  wire p1_tuple_index_1492_comb;
  wire p1_tuple_index_1493_comb;
  wire [27:0] p1_wide_x__1_comb;
  wire p1_x_sign_comb;
  wire p1_y_sign_comb;
  wire [27:0] p1_neg_1499_comb;
  wire [27:0] p1_sticky_comb;
  wire [27:0] p1_addend_y__2_comb;
  wire [24:0] p1_sel_1506_comb;
  wire [25:0] p1_add_1511_comb;
  wire [27:0] p1_concat_1514_comb;
  wire [27:0] p1_abs_fraction__2_comb;
  wire [27:0] p1_reverse_1518_comb;
  wire [28:0] p1_one_hot_1519_comb;
  wire [4:0] p1_encode_1520_comb;
  wire p1_cancel__2_comb;
  wire p1_carry_bit_comb;
  wire [27:0] p1_leading_zeroes_comb;
  wire [26:0] p1_carry_fraction_comb;
  wire [27:0] p1_add_1537_comb;
  wire [2:0] p1_concat_1538_comb;
  wire [26:0] p1_carry_fraction__1_comb;
  wire [26:0] p1_cancel_fraction_comb;
  wire [26:0] p1_shifted_fraction_comb;
  wire [2:0] p1_normal_chunk_comb;
  wire [1:0] p1_half_way_chunk_comb;
  wire [24:0] p1_add_1553_comb;
  wire p1_do_round_up_comb;
  wire [27:0] p1_rounded_fraction_comb;
  wire p1_rounding_carry_comb;
  wire [8:0] p1_add_1564_comb;
  wire [9:0] p1_add_1572_comb;
  wire [9:0] p1_wide_exponent_comb;
  wire [9:0] p1_wide_exponent__1_comb;
  wire [7:0] p1_MAX_EXPONENT__8_comb;
  wire [7:0] p1_MAX_EXPONENT__9_comb;
  wire [7:0] p1_MAX_EXPONENT__3_comb;
  wire [7:0] p1_MAX_EXPONENT__6_comb;
  wire p1_ne_1593_comb;
  wire p1_ne_1595_comb;
  wire p1_eq_1596_comb;
  wire p1_eq_1597_comb;
  wire p1_eq_1598_comb;
  wire p1_eq_1599_comb;
  wire [8:0] p1_wide_exponent__2_comb;
  wire p1_fraction_is_zero_comb;
  wire p1_has_pos_inf_comb;
  wire p1_has_neg_inf_comb;
  wire [2:0] p1_fraction_shift__1_comb;
  wire p1_and_reduce_1620_comb;
  wire p1_and_1621_comb;
  wire p1_and_1622_comb;
  wire [2:0] p1_concat_1626_comb;
  wire [27:0] p1_shrl_1629_comb;
  wire p1_is_result_nan_comb;
  wire p1_is_operand_inf_comb;
  wire p1_result_sign_comb;
  wire [22:0] p1_result_fraction_comb;
  wire p1_result_sign__1_comb;
  wire [7:0] p1_MAX_EXPONENT__7_comb;
  wire [22:0] p1_result_fraction__3_comb;
  wire [22:0] p1_FRACTION_HIGH_BIT_comb;
  wire p1_result_sign__2_comb;
  wire [7:0] p1_result_exponent__2_comb;
  wire [22:0] p1_result_fraction__4_comb;
  wire [31:0] p1_tuple_1653_comb;
  assign p1_b_bexp__2_comb = p0_b[30:23];
  assign p1_a_bexp__2_comb = p0_a[30:23];
  assign p1_sum_comb = {1'h0, p1_a_bexp__2_comb} + {1'h0, ~p1_b_bexp__2_comb};
  assign p1_tuple_index_1463_comb = p0_a[22:0];
  assign p1_tuple_index_1464_comb = p0_b[22:0];
  assign p1_y_bexp_comb = p1_sum_comb[8] ? p1_b_bexp__2_comb : p1_a_bexp__2_comb;
  assign p1_y_fraction_comb = p1_sum_comb[8] ? p1_tuple_index_1464_comb : p1_tuple_index_1463_comb;
  assign p1_incremented_sum__1_comb = p1_sum_comb[7:0] + 8'h01;
  assign p1_wide_y_comb = {2'h1, p1_y_fraction_comb, 3'h0};
  assign p1_a_bexpbs_difference__1_comb = p1_sum_comb[8] ? p1_incremented_sum__1_comb : ~p1_sum_comb[7:0];
  assign p1_x_bexp_comb = p1_sum_comb[8] ? p1_a_bexp__2_comb : p1_b_bexp__2_comb;
  assign p1_wide_y__1_comb = p1_wide_y_comb & {28{p1_y_bexp_comb != 8'h00}};
  assign p1_sub_1482_comb = 8'h1c - p1_a_bexpbs_difference__1_comb;
  assign p1_x_fraction_comb = p1_sum_comb[8] ? p1_tuple_index_1463_comb : p1_tuple_index_1464_comb;
  assign p1_dropped_comb = p1_sub_1482_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__1_comb << p1_sub_1482_comb;
  assign p1_wide_x_comb = {2'h1, p1_x_fraction_comb, 3'h0};
  assign p1_tuple_index_1492_comb = p0_b[31:31];
  assign p1_tuple_index_1493_comb = p0_a[31:31];
  assign p1_wide_x__1_comb = p1_wide_x_comb & {28{p1_x_bexp_comb != 8'h00}};
  assign p1_x_sign_comb = p1_sum_comb[8] ? p1_tuple_index_1493_comb : p1_tuple_index_1492_comb;
  assign p1_y_sign_comb = p1_sum_comb[8] ? p1_tuple_index_1492_comb : p1_tuple_index_1493_comb;
  assign p1_neg_1499_comb = -p1_wide_x__1_comb;
  assign p1_sticky_comb = {27'h000_0000, p1_dropped_comb[27:3] != 25'h000_0000};
  assign p1_addend_y__2_comb = (p1_a_bexpbs_difference__1_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__1_comb >> p1_a_bexpbs_difference__1_comb) | p1_sticky_comb;
  assign p1_sel_1506_comb = p1_x_sign_comb ^ p1_y_sign_comb ? p1_neg_1499_comb[27:3] : p1_wide_x__1_comb[27:3];
  assign p1_add_1511_comb = {{1{p1_sel_1506_comb[24]}}, p1_sel_1506_comb} + {1'h0, p1_addend_y__2_comb[27:3]};
  assign p1_concat_1514_comb = {p1_add_1511_comb[24:0], p1_addend_y__2_comb[2:0]};
  assign p1_abs_fraction__2_comb = p1_add_1511_comb[25] ? -p1_concat_1514_comb : p1_concat_1514_comb;
  assign p1_reverse_1518_comb = {p1_abs_fraction__2_comb[0], p1_abs_fraction__2_comb[1], p1_abs_fraction__2_comb[2], p1_abs_fraction__2_comb[3], p1_abs_fraction__2_comb[4], p1_abs_fraction__2_comb[5], p1_abs_fraction__2_comb[6], p1_abs_fraction__2_comb[7], p1_abs_fraction__2_comb[8], p1_abs_fraction__2_comb[9], p1_abs_fraction__2_comb[10], p1_abs_fraction__2_comb[11], p1_abs_fraction__2_comb[12], p1_abs_fraction__2_comb[13], p1_abs_fraction__2_comb[14], p1_abs_fraction__2_comb[15], p1_abs_fraction__2_comb[16], p1_abs_fraction__2_comb[17], p1_abs_fraction__2_comb[18], p1_abs_fraction__2_comb[19], p1_abs_fraction__2_comb[20], p1_abs_fraction__2_comb[21], p1_abs_fraction__2_comb[22], p1_abs_fraction__2_comb[23], p1_abs_fraction__2_comb[24], p1_abs_fraction__2_comb[25], p1_abs_fraction__2_comb[26], p1_abs_fraction__2_comb[27]};
  assign p1_one_hot_1519_comb = {p1_reverse_1518_comb[27:0] == 28'h000_0000, p1_reverse_1518_comb[27] && p1_reverse_1518_comb[26:0] == 27'h000_0000, p1_reverse_1518_comb[26] && p1_reverse_1518_comb[25:0] == 26'h000_0000, p1_reverse_1518_comb[25] && p1_reverse_1518_comb[24:0] == 25'h000_0000, p1_reverse_1518_comb[24] && p1_reverse_1518_comb[23:0] == 24'h00_0000, p1_reverse_1518_comb[23] && p1_reverse_1518_comb[22:0] == 23'h00_0000, p1_reverse_1518_comb[22] && p1_reverse_1518_comb[21:0] == 22'h00_0000, p1_reverse_1518_comb[21] && p1_reverse_1518_comb[20:0] == 21'h00_0000, p1_reverse_1518_comb[20] && p1_reverse_1518_comb[19:0] == 20'h0_0000, p1_reverse_1518_comb[19] && p1_reverse_1518_comb[18:0] == 19'h0_0000, p1_reverse_1518_comb[18] && p1_reverse_1518_comb[17:0] == 18'h0_0000, p1_reverse_1518_comb[17] && p1_reverse_1518_comb[16:0] == 17'h0_0000, p1_reverse_1518_comb[16] && p1_reverse_1518_comb[15:0] == 16'h0000, p1_reverse_1518_comb[15] && p1_reverse_1518_comb[14:0] == 15'h0000, p1_reverse_1518_comb[14] && p1_reverse_1518_comb[13:0] == 14'h0000, p1_reverse_1518_comb[13] && p1_reverse_1518_comb[12:0] == 13'h0000, p1_reverse_1518_comb[12] && p1_reverse_1518_comb[11:0] == 12'h000, p1_reverse_1518_comb[11] && p1_reverse_1518_comb[10:0] == 11'h000, p1_reverse_1518_comb[10] && p1_reverse_1518_comb[9:0] == 10'h000, p1_reverse_1518_comb[9] && p1_reverse_1518_comb[8:0] == 9'h000, p1_reverse_1518_comb[8] && p1_reverse_1518_comb[7:0] == 8'h00, p1_reverse_1518_comb[7] && p1_reverse_1518_comb[6:0] == 7'h00, p1_reverse_1518_comb[6] && p1_reverse_1518_comb[5:0] == 6'h00, p1_reverse_1518_comb[5] && p1_reverse_1518_comb[4:0] == 5'h00, p1_reverse_1518_comb[4] && p1_reverse_1518_comb[3:0] == 4'h0, p1_reverse_1518_comb[3] && p1_reverse_1518_comb[2:0] == 3'h0, p1_reverse_1518_comb[2] && p1_reverse_1518_comb[1:0] == 2'h0, p1_reverse_1518_comb[1] && !p1_reverse_1518_comb[0], p1_reverse_1518_comb[0]};
  assign p1_encode_1520_comb = {p1_one_hot_1519_comb[16] | p1_one_hot_1519_comb[17] | p1_one_hot_1519_comb[18] | p1_one_hot_1519_comb[19] | p1_one_hot_1519_comb[20] | p1_one_hot_1519_comb[21] | p1_one_hot_1519_comb[22] | p1_one_hot_1519_comb[23] | p1_one_hot_1519_comb[24] | p1_one_hot_1519_comb[25] | p1_one_hot_1519_comb[26] | p1_one_hot_1519_comb[27] | p1_one_hot_1519_comb[28], p1_one_hot_1519_comb[8] | p1_one_hot_1519_comb[9] | p1_one_hot_1519_comb[10] | p1_one_hot_1519_comb[11] | p1_one_hot_1519_comb[12] | p1_one_hot_1519_comb[13] | p1_one_hot_1519_comb[14] | p1_one_hot_1519_comb[15] | p1_one_hot_1519_comb[24] | p1_one_hot_1519_comb[25] | p1_one_hot_1519_comb[26] | p1_one_hot_1519_comb[27] | p1_one_hot_1519_comb[28], p1_one_hot_1519_comb[4] | p1_one_hot_1519_comb[5] | p1_one_hot_1519_comb[6] | p1_one_hot_1519_comb[7] | p1_one_hot_1519_comb[12] | p1_one_hot_1519_comb[13] | p1_one_hot_1519_comb[14] | p1_one_hot_1519_comb[15] | p1_one_hot_1519_comb[20] | p1_one_hot_1519_comb[21] | p1_one_hot_1519_comb[22] | p1_one_hot_1519_comb[23] | p1_one_hot_1519_comb[28], p1_one_hot_1519_comb[2] | p1_one_hot_1519_comb[3] | p1_one_hot_1519_comb[6] | p1_one_hot_1519_comb[7] | p1_one_hot_1519_comb[10] | p1_one_hot_1519_comb[11] | p1_one_hot_1519_comb[14] | p1_one_hot_1519_comb[15] | p1_one_hot_1519_comb[18] | p1_one_hot_1519_comb[19] | p1_one_hot_1519_comb[22] | p1_one_hot_1519_comb[23] | p1_one_hot_1519_comb[26] | p1_one_hot_1519_comb[27], p1_one_hot_1519_comb[1] | p1_one_hot_1519_comb[3] | p1_one_hot_1519_comb[5] | p1_one_hot_1519_comb[7] | p1_one_hot_1519_comb[9] | p1_one_hot_1519_comb[11] | p1_one_hot_1519_comb[13] | p1_one_hot_1519_comb[15] | p1_one_hot_1519_comb[17] | p1_one_hot_1519_comb[19] | p1_one_hot_1519_comb[21] | p1_one_hot_1519_comb[23] | p1_one_hot_1519_comb[25] | p1_one_hot_1519_comb[27]};
  assign p1_cancel__2_comb = |p1_encode_1520_comb[4:1];
  assign p1_carry_bit_comb = p1_abs_fraction__2_comb[27];
  assign p1_leading_zeroes_comb = {23'h00_0000, p1_encode_1520_comb};
  assign p1_carry_fraction_comb = p1_abs_fraction__2_comb[27:1];
  assign p1_add_1537_comb = p1_leading_zeroes_comb + 28'hfff_ffff;
  assign p1_concat_1538_comb = {~(p1_carry_bit_comb | p1_cancel__2_comb), ~(p1_carry_bit_comb | ~p1_cancel__2_comb), ~(~p1_carry_bit_comb | p1_cancel__2_comb)};
  assign p1_carry_fraction__1_comb = p1_carry_fraction_comb | {26'h000_0000, p1_abs_fraction__2_comb[0]};
  assign p1_cancel_fraction_comb = p1_add_1537_comb >= 28'h000_001b ? 27'h000_0000 : p1_abs_fraction__2_comb[26:0] << p1_add_1537_comb;
  assign p1_shifted_fraction_comb = p1_carry_fraction__1_comb & {27{p1_concat_1538_comb[0]}} | p1_cancel_fraction_comb & {27{p1_concat_1538_comb[1]}} | p1_abs_fraction__2_comb[26:0] & {27{p1_concat_1538_comb[2]}};
  assign p1_normal_chunk_comb = p1_shifted_fraction_comb[2:0];
  assign p1_half_way_chunk_comb = p1_shifted_fraction_comb[3:2];
  assign p1_add_1553_comb = {1'h0, p1_shifted_fraction_comb[26:3]} + 25'h000_0001;
  assign p1_do_round_up_comb = p1_normal_chunk_comb > 3'h4 | p1_half_way_chunk_comb == 2'h3;
  assign p1_rounded_fraction_comb = p1_do_round_up_comb ? {p1_add_1553_comb, p1_normal_chunk_comb} : {1'h0, p1_shifted_fraction_comb};
  assign p1_rounding_carry_comb = p1_rounded_fraction_comb[27];
  assign p1_add_1564_comb = {1'h0, p1_x_bexp_comb} + {8'h00, p1_rounding_carry_comb};
  assign p1_add_1572_comb = {1'h0, p1_add_1564_comb} + 10'h001;
  assign p1_wide_exponent_comb = p1_add_1572_comb - {5'h00, p1_encode_1520_comb};
  assign p1_wide_exponent__1_comb = p1_wide_exponent_comb & {10{p1_add_1511_comb != 26'h000_0000 | p1_addend_y__2_comb[2:0] != 3'h0}};
  assign p1_MAX_EXPONENT__8_comb = 8'hff;
  assign p1_MAX_EXPONENT__9_comb = 8'hff;
  assign p1_MAX_EXPONENT__3_comb = 8'hff;
  assign p1_MAX_EXPONENT__6_comb = 8'hff;
  assign p1_ne_1593_comb = p1_x_fraction_comb != 23'h00_0000;
  assign p1_ne_1595_comb = p1_y_fraction_comb != 23'h00_0000;
  assign p1_eq_1596_comb = p1_x_bexp_comb == p1_MAX_EXPONENT__3_comb;
  assign p1_eq_1597_comb = p1_x_fraction_comb == 23'h00_0000;
  assign p1_eq_1598_comb = p1_y_bexp_comb == p1_MAX_EXPONENT__6_comb;
  assign p1_eq_1599_comb = p1_y_fraction_comb == 23'h00_0000;
  assign p1_wide_exponent__2_comb = p1_wide_exponent__1_comb[8:0] & {9{~p1_wide_exponent__1_comb[9]}};
  assign p1_fraction_is_zero_comb = p1_add_1511_comb == 26'h000_0000 & p1_addend_y__2_comb[2:0] == 3'h0;
  assign p1_has_pos_inf_comb = ~(p1_x_bexp_comb != p1_MAX_EXPONENT__8_comb | p1_ne_1593_comb | p1_x_sign_comb) | ~(p1_y_bexp_comb != p1_MAX_EXPONENT__9_comb | p1_ne_1595_comb | p1_y_sign_comb);
  assign p1_has_neg_inf_comb = p1_eq_1596_comb & p1_eq_1597_comb & p1_x_sign_comb | p1_eq_1598_comb & p1_eq_1599_comb & p1_y_sign_comb;
  assign p1_fraction_shift__1_comb = {2'h0, p1_rounding_carry_comb} + 3'h3;
  assign p1_and_reduce_1620_comb = &p1_wide_exponent__2_comb[7:0];
  assign p1_and_1621_comb = p1_eq_1596_comb & p1_eq_1597_comb;
  assign p1_and_1622_comb = p1_eq_1598_comb & p1_eq_1599_comb;
  assign p1_concat_1626_comb = {~(p1_add_1511_comb[25] | p1_fraction_is_zero_comb), p1_add_1511_comb[25], p1_fraction_is_zero_comb};
  assign p1_shrl_1629_comb = p1_rounded_fraction_comb >> p1_fraction_shift__1_comb;
  assign p1_is_result_nan_comb = p1_eq_1596_comb & p1_ne_1593_comb | p1_eq_1598_comb & p1_ne_1595_comb | p1_has_pos_inf_comb & p1_has_neg_inf_comb;
  assign p1_is_operand_inf_comb = p1_and_1621_comb | p1_and_1622_comb;
  assign p1_result_sign_comb = p1_x_sign_comb & p1_y_sign_comb & p1_concat_1626_comb[0] | ~p1_y_sign_comb & p1_concat_1626_comb[1] | p1_y_sign_comb & p1_concat_1626_comb[2];
  assign p1_result_fraction_comb = p1_shrl_1629_comb[22:0];
  assign p1_result_sign__1_comb = p1_is_operand_inf_comb ? ~p1_has_pos_inf_comb : p1_result_sign_comb;
  assign p1_MAX_EXPONENT__7_comb = 8'hff;
  assign p1_result_fraction__3_comb = p1_result_fraction_comb & {23{(|p1_wide_exponent__2_comb[8:1]) | p1_wide_exponent__2_comb[0]}} & {23{~(p1_wide_exponent__2_comb[8] | p1_and_reduce_1620_comb)}} & {23{~(p1_and_1621_comb | p1_and_1622_comb)}};
  assign p1_FRACTION_HIGH_BIT_comb = 23'h40_0000;
  assign p1_result_sign__2_comb = ~p1_is_result_nan_comb & p1_result_sign__1_comb;
  assign p1_result_exponent__2_comb = p1_is_result_nan_comb | p1_is_operand_inf_comb | p1_wide_exponent__2_comb[8] | p1_and_reduce_1620_comb ? p1_MAX_EXPONENT__7_comb : p1_wide_exponent__2_comb[7:0];
  assign p1_result_fraction__4_comb = p1_is_result_nan_comb ? p1_FRACTION_HIGH_BIT_comb : p1_result_fraction__3_comb;
  assign p1_tuple_1653_comb = {p1_result_sign__2_comb, p1_result_exponent__2_comb, p1_result_fraction__4_comb};

  // Registers for pipe stage 1:
  reg [31:0] p1_tuple_1653;
  always_ff @ (posedge clk) begin
    p1_tuple_1653 <= p1_tuple_1653_comb;
  end
  carry_and_cancel: assert property (@(posedge clk) disable iff ($isunknown(~(p1_carry_bit_comb & p1_cancel__2_comb))) ~(p1_carry_bit_comb & p1_cancel__2_comb)) else $fatal(0, "Assertion failure via fail! @ adler32.x:2522:19-2522:66");
  assign out = p1_tuple_1653;
endmodule
